library verilog;
use verilog.vl_types.all;
entity SRFLIPFLOPUSINGCASE_vlg_vec_tst is
end SRFLIPFLOPUSINGCASE_vlg_vec_tst;
